-- comparator pentru stabilirea urmatoarei destinatii a liftului in functie de prioritatea de cautare

entity comp_decizie is
	port(n2: in bit_vector (3 downto 0);   -- etajul curent
	sus: in bit_vector (12 downto 0); 	-- cererile de urcare
	jos: in bit_vector (12 downto 0);   -- cererile de coborare
	sens_lift: in bit;		   -- sensul de deplasare al liftului
	dec: out bit_vector (12 downto 0));	 -- decizia luata (urmatoarea destinatie a liftului)
end comp_decizie;

architecture arch of comp_decizie is
begin
	process (sens_lift,n2,sus,jos)
	begin
			if sens_lift='1' then	-- daca liftul urca, se vor verifica cererile dupa cum urmeaza, in ordine: cererile de urcare de la un nivel superior, cererile de coborare de la un nivel superior,
						case n2 is 	-- cererile de urcare de la un etaj inferior etajului curent, cererile de coborare de la un etaj inferior etajului curent
									-- prioritara dintre cererile de urcare este in general cea de la etajul cel mai mic, iar pentru cele de coborare cea de la etajul cel mai mare
									-- explicatia detaliata in documentatia proiectului
							when "0000" => 
							
							if sus(0)='0' then 
							if sus(1)='0' then
							if sus(2)='0' then 
							if sus(3)='0' then			
							if sus(4)='0' then
							if sus(5)='0' then
							if sus(6)='0' then
							if sus(7)='0' then
							if sus(8)='0' then
							if sus(9)='0' then
							if sus(10)='0' then
							if sus(11)='0' then
							if sus(12)='0' then
							if jos(12)='0' then	
							if jos(11)='0' then
							if jos(10)='0' then
							if jos(9)='0' then
							if jos(8)='0' then
							if jos(7)='0' then
							if jos(6)='0' then
							if jos(5)='0' then
							if jos(4)='0' then
							if jos(3)='0' then
							if jos(2)='0' then
							if jos(1)='0' then
							if jos(0)='0' then
								dec<="0000000000000"; 	-- liftul a onorat toate cererile, deci nu se va mai deplasa, ramanand la etajul curent pana la aparitia unei noi cereri
							else dec<="0000000000001"; end if;
							else dec<="0000000000010"; end if;
							else dec<="0000000000100"; end if;
							else dec<="0000000001000"; end if;
							else dec<="0000000010000"; end if;
							else dec<="0000000100000"; end if;
							else dec<="0000001000000"; end if;
							else dec<="0000010000000"; end if;	
							else dec<="0000100000000"; end if;
							else dec<="0001000000000"; end if;
							else dec<="0010000000000"; end if;	
							else dec<="0100000000000"; end if;
							else dec<="1000000000000"; end if;
							else dec<="1000000000000"; end if;
							else dec<="0100000000000"; end if;
							else dec<="0010000000000"; end if;
							else dec<="0001000000000"; end if;
							else dec<="0000100000000"; end if;
							else dec<="0000010000000"; end if;
							else dec<="0000001000000"; end if;
							else dec<="0000000100000"; end if;
							else dec<="0000000010000"; end if;
							else dec<="0000000001000"; end if;	
							else dec<="0000000000100"; end if;	
							else dec<="0000000000010"; end if;
							else dec<="0000000000001"; end if;
							
							when "0001" => 
						
								if sus(2)='0' then 
								if sus(3)='0' then
								if sus(4)='0' then
								if sus(5)='0' then
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then
								if sus(12)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if jos(5)='0' then
								if jos(4)='0' then
								if jos(3)='0' then
								if jos(2)='0' then
								if jos(0)='0' then
								if sus(0)='0' then
									dec<="0000000000000";
								else dec<="0000000000001"; end if;
								else dec<="0000000000001"; end if;	
								else dec<="0000000000100"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if; 
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000001000"; end if;	
								else dec<="0000000000100"; end if;	
							
							when "0010" => 
						
								if sus(3)='0' then
								if sus(4)='0' then
								if sus(5)='0' then
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then	
								if sus(12)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if jos(5)='0' then
								if jos(4)='0' then
								if jos(3)='0' then
								if sus(0)='0' then
								if sus(1)='0' then
								if jos(1)='0' then
								if jos(0)='0' then
									dec<="0000000000000";
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000001000"; end if;
							
							when "0011" => 
						
								if sus(4)='0' then
								if sus(5)='0' then
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then	
								if sus(12)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if jos(5)='0' then
								if jos(4)='0' then
								if sus(0)='0' then
								if sus(1)='0' then 
								if sus(2)='0' then
								if jos(2)='0' then
								if jos(1)='0' then
								if jos(0)='0' then
									dec<="0000000000000";
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000010000"; end if;	
							
							when "0100" => 
						
								if sus(5)='0' then
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then
								if sus(12)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if jos(5)='0' then
								if sus(0)='0' then
								if sus(1)='0' then 
								if sus(2)='0' then
								if sus(3)='0' then
								if jos(3)='0' then
								if jos(2)='0' then
								if jos(1)='0' then 
								if jos(0)='0' then
									dec<="0000000000000";
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000000100000"; end if;
							
							when "0101" => 
						
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then	
								if sus(12)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if sus(0)='0' then
								if sus(1)='0' then 
								if sus(2)='0' then
								if sus(3)='0' then 
								if sus(4)='0' then
								if jos(4)='0' then
								if jos(3)='0' then
								if jos(2)='0' then
								if jos(1)='0' then
								if jos(0)='0' then
									dec<="0000000000000";
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000001000"; end if;	 
								else dec<="0000000010000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if; 
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;	
							
							when "0110" => 
						
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then
								if sus(12)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if sus(0)='0' then
								if sus(1)='0' then 
								if sus(2)='0' then
								if sus(3)='0' then 
								if sus(4)='0' then
								if sus(5)='0' then
								if jos(5)='0' then
								if jos(4)='0' then
								if jos(3)='0' then
								if jos(2)='0' then
								if jos(1)='0' then 
								if jos(0)='0' then
									dec<="0000000000000";
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000001000"; end if;	 
								else dec<="0000000010000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;	 
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
							
							when "0111" => 
									if sus(8)='0' then
									if sus(9)='0' then
									if sus(10)='0' then
									if sus(11)='0' then	
									if sus(12)='0' then
									if jos(12)='0' then	
									if jos(11)='0' then
									if jos(10)='0' then
									if jos(9)='0' then
									if jos(8)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then
									if jos(0)='0' then
										dec<="0000000000000";
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000";end if;	 
									else dec<="0000000010000";end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																														
									else dec<="0000000000001"; end if;	
									else dec<="0000100000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0010000000000"; end if;	
									else dec<="0100000000000"; end if;
									else dec<="1000000000000"; end if;	
									else dec<="1000000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0000100000000"; end if;	
							
							when "1000" => 
									if sus(9)='0' then
									if sus(10)='0' then
									if sus(11)='0' then
									if sus(12)='0' then
									if jos(12)='0' then	
									if jos(11)='0' then
									if jos(10)='0' then
									if jos(9)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then
									if jos(0)='0' then
										dec<="0000000000000";
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000";end if;	 
									else dec<="0000000010000";end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																					
									else dec<="0000000000001"; end if;	
									else dec<="0001000000000"; end if;
									else dec<="0010000000000"; end if;	
									else dec<="0100000000000"; end if;
									else dec<="1000000000000"; end if;
									else dec<="1000000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0001000000000"; end if;
							
							when "1001" => 
									if sus(10)='0' then
									if sus(11)='0' then
									if sus(12)='0' then
									if jos(12)='0' then	
									if jos(11)='0' then
									if jos(10)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if sus(8)='0' then
									if jos(8)='0' then
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then 
									if jos(0)='0' then
										dec<="0000000000000";
									else dec<="0000000000001";end if;
									else dec<="0000000000010";end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000";end if;	 
									else dec<="0000000010000";end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																				
									else dec<="0000000000001"; end if;	
									else dec<="0010000000000"; end if;	
									else dec<="0100000000000"; end if;
									else dec<="1000000000000"; end if;
									else dec<="1000000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="0010000000000"; end if;	
							
							when "1010" => 
									if sus(11)='0' then
									if sus(12)='0' then
									if jos(12)='0' then	
									if jos(11)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if sus(8)='0' then
									if sus(9)='0' then
									if jos(9)='0' then
									if jos(8)='0' then
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then 
									if jos(0)='0' then
										dec<="0000000000000";
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000"; end if;	 
									else dec<="0000000010000"; end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																														
									else dec<="0000000000001"; end if;		
									else dec<="0100000000000"; end if;
									else dec<="1000000000000"; end if;
									else dec<="1000000000000"; end if;
									else dec<="0100000000000"; end if;
							
							when "1011" =>
									if sus(12)='0' then
									if jos(12)='0' then	
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if sus(8)='0' then
									if sus(9)='0' then 
									if sus(10)='0' then
									if jos(10)='0' then
									if jos(9)='0' then
									if jos(8)='0' then
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then
									if jos(0)='0' then
										dec<="0000000000000";
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000"; end if;	 
									else dec<="0000000010000"; end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																														
									else dec<="0000000000001"; end if;		
									else dec<="1000000000000"; end if; 
									else dec<="1000000000000"; end if;
							
							when "1100" => 
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if sus(8)='0' then
									if sus(9)='0' then 
									if sus(10)='0' then
									if sus(11)='0' then
									if jos(11)='0' then
									if jos(10)='0' then
									if jos(9)='0' then
									if jos(8)='0' then
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then
									if jos(0)='0' then
										dec<="0000000000000";
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000"; end if;	 
									else dec<="0000000010000"; end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000";end if;
									else dec<="0000000000100";end if;
									else dec<="0000000000010";end if;
									else dec<="0000000000001"; end if;				
							when others => null;
							end case;
					else		 -- daca liftul coboara, se vor verifica cererile dupa cum urmeaza, in ordine: cererile de coborare de la un etaj inferior, cererile de urcare de la un etaj superior,
								 -- cererile de coborare de la un nivel superior,	cererile de urcare de la un nivel superior etajului curent
						case n2 is
							when "1100" => 
									if jos(11)='0' then
									if jos(10)='0' then
									if jos(9)='0' then
									if jos(8)='0' then
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then 
									if jos(0)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if sus(8)='0' then
									if sus(9)='0' then 
									if sus(10)='0' then
									if sus(11)='0' then
										
									
										dec<="0000000000000";
									else dec<="0100000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000001"; end if;
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000"; end if;	 
									else dec<="0000000010000"; end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0100000000000"; end if;
										
							when "1011" => 
							
									if jos(10)='0' then
									if jos(9)='0' then
									if jos(8)='0' then
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then
									if jos(0)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if sus(8)='0' then
									if sus(9)='0' then 
									if sus(10)='0' then	
									if sus(12)='0' then
									if jos(12)='0' then	
										dec<="0000000000000";
									else dec<="1000000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																														
									else dec<="0000000000001"; end if;
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000"; end if;	 
									else dec<="0000000010000"; end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="1000000000000"; end if;
									  							
							when "1010" => 
							
									if jos(9)='0' then
									if jos(8)='0' then
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then
									if jos(0)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if sus(8)='0' then
									if sus(9)='0' then
									if jos(12)='0' then	
									if jos(11)='0' then
									if sus(11)='0' then	
									if sus(12)='0' then
										dec<="0000000000000";
									else dec<="1000000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="1000000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																														
									else dec<="0000000000001"; end if;
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000"; end if;	 
									else dec<="0000000010000"; end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0001000000000"; end if;
											
									
									
										
							when "1001" => 
							
									if jos(8)='0' then
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then
									if jos(0)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if sus(8)='0' then
									if jos(12)='0' then	
									if jos(11)='0' then
									if jos(10)='0' then
									if sus(10)='0' then
									if sus(11)='0' then
									if sus(12)='0' then
										dec<="0000000000000";
									else dec<="1000000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0010000000000"; end if;	
									else dec<="0100000000000"; end if;
									else dec<="1000000000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																				
									else dec<="0000000000001"; end if;	
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000"; end if;	 
									else dec<="0000000010000"; end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
									else dec<="0000100000000"; end if;
										
									
									
										
							when "1000" => 
							
									if jos(7)='0' then
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then 
									if jos(0)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if sus(7)='0' then
									if jos(12)='0' then	
									if jos(11)='0' then
									if jos(10)='0' then
									if jos(9)='0' then 
									if sus(9)='0' then
									if sus(10)='0' then
									if sus(11)='0' then
									if sus(12)='0' then
										dec<="0000000000000";
									else dec<="1000000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0010000000000"; end if;	
									else dec<="0100000000000"; end if;
									else dec<="1000000000000"; end if;	
									else dec<="0000010000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																					
									else dec<="0000000000001"; end if;
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000"; end if;	 
									else dec<="0000000010000"; end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
									else dec<="0000010000000"; end if;
										
									
									 
										
							when "0111" => 	 
							
									if jos(6)='0' then
									if jos(5)='0' then
									if jos(4)='0' then
									if jos(3)='0' then
									if jos(2)='0' then
									if jos(1)='0' then
									if jos(0)='0' then
									if sus(0)='0' then
									if sus(1)='0' then 
									if sus(2)='0' then
									if sus(3)='0' then 
									if sus(4)='0' then
									if sus(5)='0' then
									if sus(6)='0' then
									if jos(12)='0' then	
									if jos(11)='0' then
									if jos(10)='0' then
									if jos(9)='0' then
									if jos(8)='0' then
									if sus(8)='0' then
									if sus(9)='0' then
									if sus(10)='0' then
									if sus(11)='0' then	
									if sus(12)='0' then
										dec<="0000000000000";
									else dec<="1000000000000"; end if;
									else dec<="0100000000000"; end if;
									else dec<="0010000000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0000100000000"; end if;
									else dec<="0001000000000"; end if;
									else dec<="0010000000000"; end if;	
									else dec<="0100000000000"; end if;
									else dec<="1000000000000"; end if;
									else dec<="0000001000000"; end if;  
									else dec<="0000000100000"; end if;
									else dec<="0000000010000"; end if;
									else dec<="0000000001000"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000000010"; end if;																														
									else dec<="0000000000001"; end if;
									else dec<="0000000000001"; end if;
									else dec<="0000000000010"; end if;
									else dec<="0000000000100"; end if;
									else dec<="0000000001000"; end if;	 
									else dec<="0000000010000"; end if;
									else dec<="0000000100000"; end if;
									else dec<="0000001000000"; end if;
										
										
									
										
							when "0110" => 
						
								if jos(5)='0' then
								if jos(4)='0' then
								if jos(3)='0' then
								if jos(2)='0' then
								if jos(1)='0' then
								if jos(0)='0' then
								if sus(0)='0' then
								if sus(1)='0' then 
								if sus(2)='0' then
								if sus(3)='0' then 
								if sus(4)='0' then
								if sus(5)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then
								if sus(12)='0' then
									dec<="0000000000000";
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;	 
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000001000"; end if;	 
								else dec<="0000000010000"; end if;
								else dec<="0000000100000"; end if;
								
								
								
									
									
						when "0101" => 
						
								if jos(4)='0' then
								if jos(3)='0' then
								if jos(2)='0' then
								if jos(1)='0' then
								if jos(0)='0' then
								if sus(0)='0' then
								if sus(1)='0' then 
								if sus(2)='0' then
								if sus(3)='0' then 
								if sus(4)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then
								if sus(12)='0' then
									dec<="0000000000000";
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000001000"; end if;	 
								else dec<="0000000010000"; end if;
								
								
								
									
						when "0100" => 
						
								if jos(3)='0' then
								if jos(2)='0' then
								if jos(1)='0' then
								if jos(0)='0' then
								if sus(0)='0' then
								if sus(1)='0' then 
								if sus(2)='0' then
								if sus(3)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if jos(5)='0' then
								if sus(5)='0' then
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then	
								if sus(11)='0' then
								if sus(12)='0' then
									dec<="0000000000000";
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000001000"; end if;
								
								
								 
									
									
						when "0011" => 
						
							   	if jos(2)='0' then
								if jos(1)='0' then
								if jos(0)='0' then
								if sus(0)='0' then
								if sus(1)='0' then 
								if sus(2)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if jos(5)='0' then
								if jos(4)='0' then
								if sus(4)='0' then
								if sus(5)='0' then
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then	
								if sus(12)='0' then
									dec<="0000000000000";
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000100"; end if;
								
								
								
									
									
									
						when "0010" => 
						
								if jos(1)='0' then 
								if jos(0)='0' then
								if sus(0)='0' then
								if sus(1)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if jos(5)='0' then
								if jos(4)='0' then
								if jos(3)='0' then
								if sus(3)='0' then
								if sus(4)='0' then
								if sus(5)='0' then
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then
								if sus(12)='0' then
									dec<="0000000000000";
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0000000000010"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000001"; end if;
								else dec<="0000000000010"; end if;

						when "0001" => 
								if jos(0)='0' then
								if sus(0)='0' then
								if jos(12)='0' then	
								if jos(11)='0' then
								if jos(10)='0' then
								if jos(9)='0' then
								if jos(8)='0' then
								if jos(7)='0' then
								if jos(6)='0' then
								if jos(5)='0' then
								if jos(4)='0' then
								if jos(3)='0' then
								if jos(2)='0' then
								if sus(2)='0' then 
								if sus(3)='0' then
								if sus(4)='0' then
								if sus(5)='0' then
								if sus(6)='0' then
								if sus(7)='0' then
								if sus(8)='0' then
								if sus(9)='0' then
								if sus(10)='0' then
								if sus(11)='0' then
								if sus(12)='0' then
									dec<="0000000000000";
								else dec<="1000000000000"; end if;
								else dec<="0100000000000"; end if;
								else dec<="0010000000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0000100000000"; end if;
								else dec<="0000010000000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000001000"; end if;	
								else dec<="0000000000100"; end if;
								else dec<="0000000000100"; end if;
								else dec<="0000000001000"; end if;
								else dec<="0000000010000"; end if;
								else dec<="0000000100000"; end if;
								else dec<="0000001000000"; end if;
								else dec<="0000010000000"; end if;	
								else dec<="0000100000000"; end if;
								else dec<="0001000000000"; end if;
								else dec<="0010000000000"; end if;	
								else dec<="0100000000000"; end if;
								else dec<="1000000000000"; end if;
								else dec<="0000000000001"; end if; 
								else dec<="0000000000001"; end if;
								 
									
									
									
						when "0000" => 
							
							if jos(12)='0' then	
							if jos(11)='0' then
							if jos(10)='0' then
							if jos(9)='0' then
							if jos(8)='0' then
							if jos(7)='0' then
							if jos(6)='0' then
							if jos(5)='0' then
							if jos(4)='0' then
							if jos(3)='0' then
							if jos(2)='0' then
							if jos(1)='0' then
							if sus(1)='0' then
							if sus(2)='0' then 
							if sus(3)='0' then
							if sus(4)='0' then
							if sus(5)='0' then
							if sus(6)='0' then
							if sus(7)='0' then
							if sus(8)='0' then
							if sus(9)='0' then
							if sus(10)='0' then
							if sus(11)='0' then
							if sus(12)='0' then
								dec<="0000000000000"; 
							else dec<="1000000000000"; end if;
							else dec<="0100000000000"; end if;
							else dec<="0010000000000"; end if;
							else dec<="0001000000000"; end if;
							else dec<="0000100000000"; end if;
							else dec<="0000010000000"; end if;
							else dec<="0000001000000"; end if;
							else dec<="0000000100000"; end if;	
							else dec<="0000000010000"; end if;
							else dec<="0000000001000"; end if;
							else dec<="0000000000100"; end if;	
							else dec<="0000000000010"; end if;
							else dec<="0000000000010"; end if;
							else dec<="0000000000100"; end if;
							else dec<="0000000001000"; end if;
							else dec<="0000000010000"; end if;
							else dec<="0000000100000"; end if;
							else dec<="0000001000000"; end if;
							else dec<="0000010000000"; end if;
							else dec<="0000100000000"; end if;
							else dec<="0001000000000"; end if;
							else dec<="0010000000000"; end if;	
							else dec<="0100000000000"; end if;	
							else dec<="1000000000000"; end if;
						
						when others => null;
						end case;
					end if;
			end process;
		end architecture;						